LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
LIBRARY work;

ENTITY instruction_decoder_box_tb IS
END ENTITY instruction_decoder_box_tb;

architecture TB of instruction_decoder_box_tb IS

    COMPONENT instruction_decoder_box IS
        PORT (
            DECODE :  IN  STD_LOGIC;
            EXECUTE :  IN  STD_LOGIC;
            IR :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
            INPUT :  OUT  STD_LOGIC;
            OUTPUT :  OUT  STD_LOGIC;
            LOAD :  OUT  STD_LOGIC;
            ADD :  OUT  STD_LOGIC;
            JUMPZ :  OUT  STD_LOGIC;
            JUMP :  OUT  STD_LOGIC;
            JUMPNZ :  OUT  STD_LOGIC;
            JUMPC :  OUT  STD_LOGIC;
            JUMPNC :  OUT  STD_LOGIC;
            SUB :  OUT  STD_LOGIC;
            BITAND :  OUT  STD_LOGIC
        );
    END COMPONENT;

    SIGNAL INPUT, OUTPUT,LOAD,ADD, JUMPZ, JUMP, JUMPNZ, JUMPC, JUMPNC, SUB, BITAND : STD_LOGIC;    
    signal IR :  STD_LOGIC_VECTOR(7 DOWNTO 0);         
    signal DECODE  : STD_LOGIC := '0';
    signal EXECUTE  : STD_LOGIC := '0';

begin 
TB : instruction_decoder_box PORT MAP(DECODE, EXECUTE, IR, INPUT, OUTPUT, LOAD, ADD,JUMPZ, JUMP,JUMPNZ, JUMPC, JUMPNC, SUB, BITAND );



DECODE <= NOT DECODE AFTER 100 ps;
EXECUTE <= NOT DECODE AFTER 200 ps;

IR  <="00000000", "00000000" AFTER 100 ps, "00000000" AFTER 200 ps, "00000000" AFTER 300 ps, "00000000" AFTER 400 ps --LOAD
,"01000000" AFTER 500 ps, "01000000" AFTER 600 ps, "01000000" AFTER 700 ps, "01000000" AFTER 800 ps     --ADD
,"00010000" AFTER 900 ps, "00010000" AFTER 1000 ps, "00010000" AFTER 1100 ps, "00010000" AFTER 1200 ps  --AND
,"01100000" AFTER 1300 ps, "01100000" AFTER 1400 ps, "01100000" AFTER 1500 ps, "01100000" AFTER 1600 ps --SUB
,"10100000" AFTER 1700 ps, "10100000" AFTER 1800 ps, "10100000" AFTER 1900 ps, "10100000" AFTER 2000 ps --INPUT
,"11100000" AFTER 2100 ps, "11100000" AFTER 2200 ps, "11100000" AFTER 2300 ps, "11100000" AFTER 2400 ps --OUTPUT
,"10000000" AFTER 2500 ps, "10000000" AFTER 2600 ps, "10000000" AFTER 2700 ps, "10000000" AFTER 2800 ps --JUMP U
,"10010000" AFTER 2900 ps, "10010000" AFTER 3000 ps, "10010000" AFTER 3100 ps, "10010000" AFTER 3200 ps --JUMP Z
,"10011000" AFTER 3300 ps, "10011000" AFTER 3400 ps, "10011000" AFTER 3500 ps, "10011000" AFTER 3600 ps --JUMP C
,"10010100" AFTER 3700 ps, "10010100" AFTER 3800 ps, "10010100" AFTER 3900 ps, "10010100" AFTER 4000 ps --JUMP NZ
,"10011100" AFTER 4100 ps, "10011100" AFTER 4200 ps, "10011100" AFTER 4300 ps, "10011100" AFTER 4400 ps; --JUMP NC

end TB;
