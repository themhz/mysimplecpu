-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"
-- CREATED		"Mon Jan 10 00:35:41 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY instruction_decoder_v2 IS 
	PORT
	(
		A :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		INPUT :  OUT  STD_LOGIC;
		OUTPUT :  OUT  STD_LOGIC;
		LOAD :  OUT  STD_LOGIC;
		ADD :  OUT  STD_LOGIC;
		JUMP :  OUT  STD_LOGIC;
		SUB :  OUT  STD_LOGIC;
		BITAND :  OUT  STD_LOGIC;
		JUMPZ :  OUT  STD_LOGIC;
		JUMPNZ :  OUT  STD_LOGIC;
		JUMPC :  OUT  STD_LOGIC;
		JUMPNC :  OUT  STD_LOGIC;
		BITOR :  OUT  STD_LOGIC
	);
END instruction_decoder_v2;

ARCHITECTURE bdf_type OF instruction_decoder_v2 IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;


BEGIN 



INPUT <= A(7) AND SYNTHESIZED_WIRE_0 AND A(5) AND SYNTHESIZED_WIRE_1;


OUTPUT <= A(7) AND A(6) AND A(5) AND SYNTHESIZED_WIRE_2;


SYNTHESIZED_WIRE_2 <= NOT(A(4));



SYNTHESIZED_WIRE_3 <= NOT(A(7));



SYNTHESIZED_WIRE_4 <= NOT(A(6));



SYNTHESIZED_WIRE_5 <= NOT(A(5));



SYNTHESIZED_WIRE_6 <= NOT(A(4));



SYNTHESIZED_WIRE_12 <= NOT(A(7));



SYNTHESIZED_WIRE_13 <= NOT(A(5));



SYNTHESIZED_WIRE_14 <= NOT(A(4));



SYNTHESIZED_WIRE_20 <= NOT(A(6));



SYNTHESIZED_WIRE_21 <= NOT(A(5));



LOAD <= SYNTHESIZED_WIRE_3 AND SYNTHESIZED_WIRE_4 AND SYNTHESIZED_WIRE_5 AND SYNTHESIZED_WIRE_6;


SYNTHESIZED_WIRE_22 <= NOT(A(4));



SYNTHESIZED_WIRE_23 <= NOT(A(6));



SYNTHESIZED_WIRE_24 <= NOT(A(5));



SYNTHESIZED_WIRE_25 <= NOT(A(7));



SYNTHESIZED_WIRE_26 <= NOT(A(4));



SYNTHESIZED_WIRE_27 <= NOT(A(7));



SYNTHESIZED_WIRE_28 <= NOT(A(6));



SYNTHESIZED_WIRE_29 <= NOT(A(5));



JUMPZ <= SYNTHESIZED_WIRE_30 AND SYNTHESIZED_WIRE_8 AND SYNTHESIZED_WIRE_9;


JUMPNZ <= SYNTHESIZED_WIRE_30 AND SYNTHESIZED_WIRE_11 AND A(2);


ADD <= SYNTHESIZED_WIRE_12 AND A(6) AND SYNTHESIZED_WIRE_13 AND SYNTHESIZED_WIRE_14;


JUMPC <= SYNTHESIZED_WIRE_30 AND A(3) AND SYNTHESIZED_WIRE_16;


JUMPNC <= SYNTHESIZED_WIRE_30 AND A(3) AND A(2);


BITOR <= SYNTHESIZED_WIRE_18 AND A(6) AND SYNTHESIZED_WIRE_19 AND A(4);


SYNTHESIZED_WIRE_8 <= NOT(A(3));



SYNTHESIZED_WIRE_9 <= NOT(A(2));



SYNTHESIZED_WIRE_11 <= NOT(A(3));



SYNTHESIZED_WIRE_16 <= NOT(A(2));



SYNTHESIZED_WIRE_18 <= NOT(A(7));



SYNTHESIZED_WIRE_19 <= NOT(A(5));



JUMP <= A(7) AND SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_21 AND SYNTHESIZED_WIRE_22;


SYNTHESIZED_WIRE_30 <= A(7) AND SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_24 AND A(4);


SUB <= SYNTHESIZED_WIRE_25 AND A(6) AND A(5) AND SYNTHESIZED_WIRE_26;


BITAND <= SYNTHESIZED_WIRE_27 AND SYNTHESIZED_WIRE_28 AND SYNTHESIZED_WIRE_29 AND A(4);


SYNTHESIZED_WIRE_0 <= NOT(A(6));



SYNTHESIZED_WIRE_1 <= NOT(A(4));



END bdf_type;