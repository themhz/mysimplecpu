-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"
-- CREATED		"Mon Jan 10 01:20:39 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY decoder_v2 IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		CE :  IN  STD_LOGIC;
		CLR :  IN  STD_LOGIC;
		Carry :  IN  STD_LOGIC;
		Zero :  IN  STD_LOGIC;
		IR :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		EN_IN :  OUT  STD_LOGIC;
		RAM :  OUT  STD_LOGIC;
		ALU_S2 :  OUT  STD_LOGIC;
		ALU_S4 :  OUT  STD_LOGIC;
		MUXA :  OUT  STD_LOGIC;
		MUXC :  OUT  STD_LOGIC;
		ALU_S1 :  OUT  STD_LOGIC;
		ALU_S0 :  OUT  STD_LOGIC;
		MUXB :  OUT  STD_LOGIC;
		EN_PC :  OUT  STD_LOGIC;
		ALU_S3 :  OUT  STD_LOGIC;
		EN_DA :  OUT  STD_LOGIC;
		ALU_S5 :  OUT  STD_LOGIC
	);
END decoder_v2;

ARCHITECTURE bdf_type OF decoder_v2 IS 

COMPONENT instruction_decoder_box_v2
	PORT(DECODE : IN STD_LOGIC;
		 EXECUTE : IN STD_LOGIC;
		 IR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 INPUT : OUT STD_LOGIC;
		 OUTPUT : OUT STD_LOGIC;
		 LOAD : OUT STD_LOGIC;
		 ADD : OUT STD_LOGIC;
		 JUMPZ : OUT STD_LOGIC;
		 JUMP : OUT STD_LOGIC;
		 JUMPNZ : OUT STD_LOGIC;
		 JUMPC : OUT STD_LOGIC;
		 JUMPNC : OUT STD_LOGIC;
		 SUB : OUT STD_LOGIC;
		 BITAND : OUT STD_LOGIC;
		 BITOR : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT status_register_v2
	PORT(Carry : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 Zero : IN STD_LOGIC;
		 ADD : IN STD_LOGIC;
		 SUB : IN STD_LOGIC;
		 BITAND : IN STD_LOGIC;
		 BITOR : IN STD_LOGIC;
		 CARRY_REG : OUT STD_LOGIC;
		 ZERO_REG : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT jump_detector
	PORT(INCREMENT : IN STD_LOGIC;
		 EXECUTE : IN STD_LOGIC;
		 ZERO_REG : IN STD_LOGIC;
		 CARRY_REG : IN STD_LOGIC;
		 JUMPZ : IN STD_LOGIC;
		 JUMPNZ : IN STD_LOGIC;
		 JUMPC : IN STD_LOGIC;
		 JUMPNC : IN STD_LOGIC;
		 JUMP : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 EN_PC : OUT STD_LOGIC;
		 jump_not_taken : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT sequence_generator
	PORT(CLK : IN STD_LOGIC;
		 CE : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 FETCH : OUT STD_LOGIC;
		 DECODE : OUT STD_LOGIC;
		 EXECUTE : OUT STD_LOGIC;
		 INCREMENT : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_13 <= '0';
SYNTHESIZED_WIRE_78 <= '0';



SYNTHESIZED_WIRE_59 <= SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64;


b2v_inst1 : instruction_decoder_box_v2
PORT MAP(DECODE => SYNTHESIZED_WIRE_2,
		 EXECUTE => SYNTHESIZED_WIRE_63,
		 IR => IR,
		 INPUT => SYNTHESIZED_WIRE_72,
		 OUTPUT => SYNTHESIZED_WIRE_64,
		 LOAD => SYNTHESIZED_WIRE_74,
		 ADD => SYNTHESIZED_WIRE_76,
		 JUMPZ => SYNTHESIZED_WIRE_67,
		 JUMP => SYNTHESIZED_WIRE_71,
		 JUMPNZ => SYNTHESIZED_WIRE_69,
		 JUMPC => SYNTHESIZED_WIRE_68,
		 JUMPNC => SYNTHESIZED_WIRE_70,
		 SUB => SYNTHESIZED_WIRE_65,
		 BITAND => SYNTHESIZED_WIRE_75,
		 BITOR => SYNTHESIZED_WIRE_77);


SYNTHESIZED_WIRE_60 <= SYNTHESIZED_WIRE_65 OR SYNTHESIZED_WIRE_66;

ALU_S4 <= SYNTHESIZED_WIRE_66;


MUXA <= SYNTHESIZED_WIRE_66;



SYNTHESIZED_WIRE_73 <= SYNTHESIZED_WIRE_67 OR SYNTHESIZED_WIRE_68 OR SYNTHESIZED_WIRE_69 OR SYNTHESIZED_WIRE_70 OR SYNTHESIZED_WIRE_71 OR SYNTHESIZED_WIRE_13;


SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_64 OR SYNTHESIZED_WIRE_72;

MUXC <= SYNTHESIZED_WIRE_16;


ALU_S1 <= SYNTHESIZED_WIRE_17;



SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_73 OR SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_75 OR SYNTHESIZED_WIRE_72;

ALU_S0 <= SYNTHESIZED_WIRE_22;



SYNTHESIZED_WIRE_17 <= SYNTHESIZED_WIRE_73 OR SYNTHESIZED_WIRE_64 OR SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_72;

MUXB <= SYNTHESIZED_WIRE_27;



b2v_inst2 : status_register_v2
PORT MAP(Carry => Carry,
		 CLK => CLK,
		 CLR => CLR,
		 Zero => Zero,
		 ADD => SYNTHESIZED_WIRE_76,
		 SUB => SYNTHESIZED_WIRE_65,
		 BITAND => SYNTHESIZED_WIRE_75,
		 BITOR => SYNTHESIZED_WIRE_77,
		 CARRY_REG => SYNTHESIZED_WIRE_51,
		 ZERO_REG => SYNTHESIZED_WIRE_50);


ALU_S3 <= SYNTHESIZED_WIRE_65;


ALU_S5 <= SYNTHESIZED_WIRE_77;



SYNTHESIZED_WIRE_27 <= SYNTHESIZED_WIRE_78 OR SYNTHESIZED_WIRE_76 OR SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_65 OR SYNTHESIZED_WIRE_75 OR SYNTHESIZED_WIRE_77;


SYNTHESIZED_WIRE_62 <= SYNTHESIZED_WIRE_78 OR SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_72 OR SYNTHESIZED_WIRE_76 OR SYNTHESIZED_WIRE_75 OR SYNTHESIZED_WIRE_65 OR SYNTHESIZED_WIRE_77 OR SYNTHESIZED_WIRE_78;


b2v_inst4 : jump_detector
PORT MAP(INCREMENT => SYNTHESIZED_WIRE_66,
		 EXECUTE => SYNTHESIZED_WIRE_63,
		 ZERO_REG => SYNTHESIZED_WIRE_50,
		 CARRY_REG => SYNTHESIZED_WIRE_51,
		 JUMPZ => SYNTHESIZED_WIRE_67,
		 JUMPNZ => SYNTHESIZED_WIRE_69,
		 JUMPC => SYNTHESIZED_WIRE_68,
		 JUMPNC => SYNTHESIZED_WIRE_70,
		 JUMP => SYNTHESIZED_WIRE_71,
		 CLK => CLK,
		 CLR => CLR,
		 EN_PC => EN_PC);


EN_IN <= SYNTHESIZED_WIRE_57;


EN_DA <= SYNTHESIZED_WIRE_58;


RAM <= SYNTHESIZED_WIRE_59;


ALU_S2 <= SYNTHESIZED_WIRE_60;



b2v_inst_sg : sequence_generator
PORT MAP(CLK => CLK,
		 CE => CE,
		 CLR => CLR,
		 FETCH => SYNTHESIZED_WIRE_57,
		 DECODE => SYNTHESIZED_WIRE_2,
		 EXECUTE => SYNTHESIZED_WIRE_63,
		 INCREMENT => SYNTHESIZED_WIRE_66);


SYNTHESIZED_WIRE_58 <= SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_62;


END bdf_type;