Library IEEE;
Use IEEE.std_logic_1164.all;
Use IEEE.std_logic_unsigned.all;

Entity RAM is
Port(din: In std_logic_vector (15 downto 0);
    addr: In std_logic_vector (7 downto 0);
    we, clk : In std_logic;
    dout: Out std_logic_vector (15 downto 0));
End RAM;

Architecture mem256x16_v2_rtl of RAM is

Type vector_array is array (0 to 255) of std_logic_vector (15 downto 0);

-- signal memory : vector_array:=(
--     0=> "1010000000001010",
--     1=> "0100000000001010",
--     2=> "1001110000000100",
--     3=> "0000000011111111",
--     4=> "1110000000001010",
--     5=> "1000000000000000",
--     6=> "0000000000000000",
--     7=> "0000000000000000",
--     8=> "0000000000000000",
--     9=> "0000000000000000",
--     10=> "0000000010000000",
--     others => "0000000000000000");

-- signal memory : vector_array:=(
--     0=> "0000000000000010",
--     1=> "0100000000000001",
--     2=> "0100000000000001",
--     others=> "0000000000000000");

-- signal memory : vector_array:=(
--     0=> "0000000000000001",
--     1=> "0100000010000001",
--     2=> "1001110000000001",
--     3=> "0000000000000000",
--     4=> "0000000000000000",
--     5=> "0000000000000000",
--     others=> "0000000000000000");

-- signal memory : vector_array:=(others=> "0000000000000000");
-- signal memory : vector_array:=(
--     0=> "0000000000110101",
--     1=> "0101000010000000",
--     others=> "0000000000000000");

-- signal memory : vector_array:=(
--     0=> "1010000001100100", --Input ACC, A064
--     1=> "0100000000000010", --Add ACC, 02
--     2=> "1110000001111001", --Output ACC,
--     3=> "1001110000000001",
--     4=> "1010000010010111",
--     5=> "1110000010010101",
--     6=> "1000000000000000",
--     151=> "0000000001001011",
--     100=> "0000000011101001",
--     others => "0000000000000000");

-- signal memory : vector_array:=(
--     0 => "0000000000000001", --LOAD ACC, 01
--     --1 => "0100000000000000", --ADD ACC, 00 // test NZ NC ACC=01
--     1 => "0100000011111111", --ADD ACC, 00 // test NZ NC ACC=01
--     2 => "1001010000001010", --JUMP NZ, 10 // skip trap if correct
--     3 => "1001000000001111", --JUMP Z, F // skip trap if correct
--     10=> "0000000000001010",
--     15=> "0000000000001101",
--     others => "0000000000000000");


-- signal memory : vector_array:=(
--     0 => "0000000010100101", --LOAD ACC, 165
--     1 => "0001000000000101", --
--     others => "0000000000000000");

signal memory : vector_array:=(
    0 => "0000000000000001", --LOAD ACC, 01
    1 => "0100000000000000", --ADD ACC, 00
    2 => "0100000011111111",--ADD ACC, FF
    3 => "0000000010101010",--LOAD ACC, AA
    4 => "0001000000001111",--AND ACC, 0F
    5 => "0001000000000000",--AND ACC, 00
    6 => "0000000000000001", --LOAD ACC, 01
    7 => "0110000000000001", --SUB ACC, 01
    8 => "0110000000000001", --SUB ACC, 01
    9 => "1001000011110000", --OUTPUT ACC, F0
    10 => "0000000000000000", --LOAD ACC, 00
    11 => "1010000011111111", --INPUT ACC, FF
    12 => "0100000000000001", --ADD ACC, 00
    13 => "1001010000001111", --JUMP NZ, 0F
    14 => "1000000000001110", --JUMP 0E
    15 => "0100000000000001", --ADD ACC, 01
    16 => "1001000000010010", --JUMP Z, 12
    17 => "1001000000010001", --JUMP NZ, 0F
    18 => "0000000000000010", --LOAD ACC, 02
    19 => "0100000011111111", --ADD ACC, FF
    20 => "1001100000010110", --JUMP C, 16
    21 => "1000000000010101", --JUMP 15
    22 => "0110000000000001", --SUB ACC, 01
    23 => "1001110000011001", --JUMP NC, 19
    24 => "1000000000011000", --TRAP
    25 => "1000000000000000", --JUMP 00    
    240 => "0000000011111111", 
    others => "0000000000000000");


    -- memory(151) <= "0000000001001011";
    -- memory(100) <= "0000000011101001";
Begin
Process (clk)
Begin
IF rising_edge(clk) then
    IF (we = '1') then
        memory(conv_integer(addr)) <= din;
    End IF;
End IF;
End Process;

dout <= memory(conv_integer(addr));

End mem256x16_v2_rtl;

