-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"
-- CREATED		"Tue Jan 04 03:19:36 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY decoder IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		CE :  IN  STD_LOGIC;
		CLR :  IN  STD_LOGIC;
		Carry :  IN  STD_LOGIC;
		Zero :  IN  STD_LOGIC;
		IR :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		EN_IN :  OUT  STD_LOGIC;
		RAM :  OUT  STD_LOGIC;
		ALU_S2 :  OUT  STD_LOGIC;
		ALU_S4 :  OUT  STD_LOGIC;
		MUXA :  OUT  STD_LOGIC;
		MUXC :  OUT  STD_LOGIC;
		ALU_S1 :  OUT  STD_LOGIC;
		ALU_S0 :  OUT  STD_LOGIC;
		MUXB :  OUT  STD_LOGIC;
		EN_PC :  OUT  STD_LOGIC;
		ALU_S3 :  OUT  STD_LOGIC;
		EN_DA :  OUT  STD_LOGIC
	);
END decoder;

ARCHITECTURE bdf_type OF decoder IS 

COMPONENT status_register
	PORT(Carry : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 Zero : IN STD_LOGIC;
		 ADD : IN STD_LOGIC;
		 SUB : IN STD_LOGIC;
		 BITAND : IN STD_LOGIC;
		 CARRY_REG : OUT STD_LOGIC;
		 ZERO_REG : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT instruction_decoder_box
	PORT(DECODE : IN STD_LOGIC;
		 EXECUTE : IN STD_LOGIC;
		 IR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 INPUT : OUT STD_LOGIC;
		 OUTPUT : OUT STD_LOGIC;
		 LOAD : OUT STD_LOGIC;
		 ADD : OUT STD_LOGIC;
		 JUMPZ : OUT STD_LOGIC;
		 JUMP : OUT STD_LOGIC;
		 JUMPNZ : OUT STD_LOGIC;
		 JUMPC : OUT STD_LOGIC;
		 JUMPNC : OUT STD_LOGIC;
		 SUB : OUT STD_LOGIC;
		 BITAND : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT jump_detector
	PORT(INCREMENT : IN STD_LOGIC;
		 EXECUTE : IN STD_LOGIC;
		 ZERO_REG : IN STD_LOGIC;
		 CARRY_REG : IN STD_LOGIC;
		 JUMPZ : IN STD_LOGIC;
		 JUMPNZ : IN STD_LOGIC;
		 JUMPC : IN STD_LOGIC;
		 JUMPNC : IN STD_LOGIC;
		 JUMP : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 EN_PC : OUT STD_LOGIC;
		 jump_not_taken : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT sequence_generator
	PORT(CLK : IN STD_LOGIC;
		 CE : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 FETCH : OUT STD_LOGIC;
		 DECODE : OUT STD_LOGIC;
		 EXECUTE : OUT STD_LOGIC;
		 INCREMENT : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_11 <= '0';
SYNTHESIZED_WIRE_17 <= '0';



SYNTHESIZED_WIRE_53 <= SYNTHESIZED_WIRE_57 AND SYNTHESIZED_WIRE_58;


SYNTHESIZED_WIRE_54 <= SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_60;

ALU_S4 <= SYNTHESIZED_WIRE_60;


MUXA <= SYNTHESIZED_WIRE_60;



SYNTHESIZED_WIRE_70 <= SYNTHESIZED_WIRE_61 OR SYNTHESIZED_WIRE_62 OR SYNTHESIZED_WIRE_63 OR SYNTHESIZED_WIRE_64 OR SYNTHESIZED_WIRE_65 OR SYNTHESIZED_WIRE_11;


SYNTHESIZED_WIRE_56 <= SYNTHESIZED_WIRE_66 OR SYNTHESIZED_WIRE_67 OR SYNTHESIZED_WIRE_68 OR SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_69 OR SYNTHESIZED_WIRE_17;


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_58 OR SYNTHESIZED_WIRE_66;

MUXC <= SYNTHESIZED_WIRE_20;


ALU_S1 <= SYNTHESIZED_WIRE_21;



SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_70 OR SYNTHESIZED_WIRE_68 OR SYNTHESIZED_WIRE_69 OR SYNTHESIZED_WIRE_66;

ALU_S0 <= SYNTHESIZED_WIRE_26;



SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_70 OR SYNTHESIZED_WIRE_58 OR SYNTHESIZED_WIRE_58 OR SYNTHESIZED_WIRE_66;

MUXB <= SYNTHESIZED_WIRE_31;



b2v_inst2 : status_register
PORT MAP(Carry => Carry,
		 CLK => CLK,
		 CLR => CLR,
		 Zero => Zero,
		 ADD => SYNTHESIZED_WIRE_67,
		 SUB => SYNTHESIZED_WIRE_59,
		 BITAND => SYNTHESIZED_WIRE_69,
		 CARRY_REG => SYNTHESIZED_WIRE_45,
		 ZERO_REG => SYNTHESIZED_WIRE_44);



SYNTHESIZED_WIRE_31 <= SYNTHESIZED_WIRE_68 OR SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_69 OR SYNTHESIZED_WIRE_67;

ALU_S3 <= SYNTHESIZED_WIRE_59;



b2v_inst3 : instruction_decoder_box
PORT MAP(DECODE => SYNTHESIZED_WIRE_40,
		 EXECUTE => SYNTHESIZED_WIRE_57,
		 IR => IR,
		 INPUT => SYNTHESIZED_WIRE_66,
		 OUTPUT => SYNTHESIZED_WIRE_58,
		 LOAD => SYNTHESIZED_WIRE_68,
		 ADD => SYNTHESIZED_WIRE_67,
		 JUMPZ => SYNTHESIZED_WIRE_61,
		 JUMP => SYNTHESIZED_WIRE_65,
		 JUMPNZ => SYNTHESIZED_WIRE_63,
		 JUMPC => SYNTHESIZED_WIRE_62,
		 JUMPNC => SYNTHESIZED_WIRE_64,
		 SUB => SYNTHESIZED_WIRE_59,
		 BITAND => SYNTHESIZED_WIRE_69);


b2v_inst4 : jump_detector
PORT MAP(INCREMENT => SYNTHESIZED_WIRE_60,
		 EXECUTE => SYNTHESIZED_WIRE_57,
		 ZERO_REG => SYNTHESIZED_WIRE_44,
		 CARRY_REG => SYNTHESIZED_WIRE_45,
		 JUMPZ => SYNTHESIZED_WIRE_61,
		 JUMPNZ => SYNTHESIZED_WIRE_63,
		 JUMPC => SYNTHESIZED_WIRE_62,
		 JUMPNC => SYNTHESIZED_WIRE_64,
		 JUMP => SYNTHESIZED_WIRE_65,
		 CLK => CLK,
		 CLR => CLR,
		 EN_PC => EN_PC);


EN_IN <= SYNTHESIZED_WIRE_51;


EN_DA <= SYNTHESIZED_WIRE_52;


RAM <= SYNTHESIZED_WIRE_53;


ALU_S2 <= SYNTHESIZED_WIRE_54;



b2v_inst_sg : sequence_generator
PORT MAP(CLK => CLK,
		 CE => CE,
		 CLR => CLR,
		 FETCH => SYNTHESIZED_WIRE_51,
		 DECODE => SYNTHESIZED_WIRE_40,
		 EXECUTE => SYNTHESIZED_WIRE_57,
		 INCREMENT => SYNTHESIZED_WIRE_60);


SYNTHESIZED_WIRE_52 <= SYNTHESIZED_WIRE_57 AND SYNTHESIZED_WIRE_56;


END bdf_type;